* File: hw2_XOR.pex.cir
* Created: Fri Nov 15 23:33:33 2024
* Program "Calibre xRC"
* Version "v2020.2_14.12"
* 
.include "hw2_XOR.pex.cir.pex"
.subckt HW2_XOR  A B C S GND VDD
* 
* VDD	VDD
* GND	GND
* S	S
* C	C
* B	B
* A	A
M0 N_5_M0_d N_B_M0_g N_3_M0_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.35e-13
+ AS=2.35e-13 PD=1.47e-06 PS=1.47e-06
M1 N_GND_M1_d N_A_M1_g N_7_M1_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.222e-13
+ AS=2.397e-13 PD=5.2e-07 PS=1.49e-06
M2 N_3_M2_d N_A_M2_g N_GND_M2_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.222e-13 PD=5.1e-07 PS=5.2e-07
M3 N_9_M3_d N_8_M3_g N_3_M3_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.2925e-13
+ AS=1.1985e-13 PD=5.5e-07 PS=5.1e-07
M4 N_S_M4_d N_C_M4_g N_9_M4_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13
+ AS=1.2925e-13 PD=5.1e-07 PS=5.5e-07
M5 N_5_M5_d N_13_M5_g N_S_M5_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.2455e-13
+ AS=1.1985e-13 PD=5.3e-07 PS=5.1e-07
M6 N_14_M6_d N_8_M6_g N_5_M6_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13
+ AS=1.2455e-13 PD=5.4e-07 PS=5.3e-07
M7 N_GND_M7_d N_7_M7_g N_14_M7_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
M8 N_14_M8_d N_B_M8_g N_9_M8_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
M9 N_GND_M9_d N_B_M9_g N_8_M9_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13
+ AS=2.303e-13 PD=5.4e-07 PS=1.45e-06
M10 N_13_M10_d N_C_M10_g N_GND_M10_s N_GND_M0_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.35e-13 AS=1.269e-13 PD=1.47e-06 PS=5.4e-07
M11 N_6_M11_d N_B_M11_g N_4_M11_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.35e-13 AS=2.35e-13 PD=1.47e-06 PS=1.47e-06
M12 N_VDD_M12_d N_A_M12_g N_7_M12_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.222e-13 AS=2.397e-13 PD=5.2e-07 PS=1.49e-06
M13 N_4_M13_d N_A_M13_g N_VDD_M13_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.222e-13 PD=5.1e-07 PS=5.2e-07
M14 N_10_M14_d N_8_M14_g N_4_M14_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.2925e-13 AS=1.1985e-13 PD=5.5e-07 PS=5.1e-07
M15 N_S_M15_d N_C_M15_g N_10_M15_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.2925e-13 PD=5.1e-07 PS=5.5e-07
M16 N_6_M16_d N_13_M16_g N_S_M16_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.2455e-13 AS=1.1985e-13 PD=5.3e-07 PS=5.1e-07
M17 N_15_M17_d N_8_M17_g N_6_M17_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=1.2455e-13 PD=5.4e-07 PS=5.3e-07
M18 N_VDD_M18_d N_7_M18_g N_15_M18_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.269e-13 PD=1.45e-06 PS=5.4e-07
M19 N_15_M19_d N_B_M19_g N_10_M19_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
M20 N_VDD_M20_d N_B_M20_g N_8_M20_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.269e-13 AS=2.303e-13 PD=5.4e-07 PS=1.45e-06
M21 N_13_M21_d N_C_M21_g N_VDD_M21_s N_VDD_M11_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.35e-13 AS=1.269e-13 PD=1.47e-06 PS=5.4e-07
*
.include "hw2_XOR.pex.cir.HW2_XOR.pxi"
*
.ends
*
*
