* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT 3XOR
** N=11 EP=0 IP=0 FDC=22
M0 5 2 3 7 N_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=2.35e-13 PD=1.02e-06 PS=1.47e-06 $X=-9780 $Y=-1390 $D=0
M1 7 1 5 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.222e-13 AS=2.397e-13 PD=5.2e-07 PS=1.02e-06 $X=-8580 $Y=-1390 $D=0
M2 3 1 7 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.222e-13 PD=5.1e-07 PS=5.2e-07 $X=-7880 $Y=-1390 $D=0
M3 7 6 3 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.2925e-13 AS=1.1985e-13 PD=5.5e-07 PS=5.1e-07 $X=-7190 $Y=-1390 $D=0
M4 10 9 7 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.2925e-13 PD=5.1e-07 PS=5.5e-07 $X=-6460 $Y=-1390 $D=0
M5 5 11 10 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.2455e-13 AS=1.1985e-13 PD=5.3e-07 PS=5.1e-07 $X=-5770 $Y=-1390 $D=0
M6 6 6 5 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.2455e-13 PD=5.4e-07 PS=5.3e-07 $X=-5060 $Y=-1390 $D=0
M7 7 5 6 7 N_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=1.269e-13 PD=9.9e-07 PS=5.4e-07 $X=-4340 $Y=-1390 $D=0
M8 6 2 7 7 N_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=2.3265e-13 PD=9.9e-07 PS=9.9e-07 $X=-3170 $Y=-1390 $D=0
M9 7 2 6 7 N_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.3265e-13 PD=5.4e-07 PS=9.9e-07 $X=-2000 $Y=-1390 $D=0
M10 11 9 7 7 N_18 L=1.8e-07 W=4.7e-07 AD=4.23e-13 AS=1.269e-13 PD=2.27e-06 PS=5.4e-07 $X=-1280 $Y=-1390 $D=0
M11 5 2 4 8 P_18 L=1.8e-07 W=4.7e-07 AD=2.397e-13 AS=2.35e-13 PD=1.02e-06 PS=1.47e-06 $X=-9780 $Y=4350 $D=1
M12 8 1 5 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.222e-13 AS=2.397e-13 PD=5.2e-07 PS=1.02e-06 $X=-8580 $Y=4350 $D=1
M13 4 1 8 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.222e-13 PD=5.1e-07 PS=5.2e-07 $X=-7880 $Y=4350 $D=1
M14 8 6 4 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.2925e-13 AS=1.1985e-13 PD=5.5e-07 PS=5.1e-07 $X=-7190 $Y=4350 $D=1
M15 10 9 8 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.1985e-13 AS=1.2925e-13 PD=5.1e-07 PS=5.5e-07 $X=-6460 $Y=4350 $D=1
M16 5 11 10 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.2455e-13 AS=1.1985e-13 PD=5.3e-07 PS=5.1e-07 $X=-5770 $Y=4350 $D=1
M17 6 6 5 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=1.2455e-13 PD=5.4e-07 PS=5.3e-07 $X=-5060 $Y=4350 $D=1
M18 8 5 6 8 P_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=1.269e-13 PD=9.9e-07 PS=5.4e-07 $X=-4340 $Y=4350 $D=1
M19 6 2 8 8 P_18 L=1.8e-07 W=4.7e-07 AD=2.3265e-13 AS=2.3265e-13 PD=9.9e-07 PS=9.9e-07 $X=-3170 $Y=4350 $D=1
M20 8 2 6 8 P_18 L=1.8e-07 W=4.7e-07 AD=1.269e-13 AS=2.3265e-13 PD=5.4e-07 PS=9.9e-07 $X=-2000 $Y=4350 $D=1
M21 11 9 8 8 P_18 L=1.8e-07 W=4.7e-07 AD=4.23e-13 AS=1.269e-13 PD=2.27e-06 PS=5.4e-07 $X=-1280 $Y=4350 $D=1
.ENDS
***************************************
